-- Instruction-Level Power Side-Channel Leakage Evaluation of Soft-Core CPUs on Shared FPGAs
-- Copyright 2023, School of Computer and Communication Sciences, EPFL.
--
-- All rights reserved. Use of this source code is governed by a
-- BSD-style license that can be found in the LICENSE.md file.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CPU_tb is
--  Port ( );
end CPU_tb;

architecture Behavioral of CPU_tb is

signal Kin, Din : std_logic_vector(127 downto 0);
signal clk, reset_n, Drdy, krdy, sensor_fifo_read, bsy, en_cpu: std_logic;
signal kvld, sensor_trigger, calib_trg, fsm_dvld, dvld_mux, rst_cpu, reset_fifo, sensor_fifo_dvld, osc_trigger: std_logic;
signal instruction_processed : std_logic_vector(31 downto 0);
signal sens_calib_id : std_logic_vector(4 downto 0);

type sig_array_lw_add is array (1 to 16) of std_logic_vector(127 downto 0);
signal instrs_lw_add : sig_array_lw_add := (
X"0000253700c54513038485b700000000",
X"0d45c593cd136db782fdcd9300000001",
X"041841b71001c1930c1ecc3700000001",
X"1a9c4c1300003d37ffbd4d1300000001",
X"00080e37ff7e4e130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00052e0301ac01b303b5d46300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e000000130000001300000001",
X"0000007e0000007e0000007efffffff2"
);

type sig_array_sw_add is array (1 to 13) of std_logic_vector(127 downto 0);
signal instrs_sw_add : sig_array_sw_add := (
X"ffff7737b8c7471348f8113700000000",
X"b8414113048803370213431300000001",
X"c2c843b71cf3c39301000ab700000001",
X"ffbaca9350ce2db7f97dcd9300000001",
X"086c0eb7fffece9301004f3700000001",
X"ffff4f13000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"01e7202301d303b341bad13300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e000000130000001300000001",
X"0000007e0000007e0000007efffffff2"
);

type sig_array is array (1 to 19) of std_logic_vector(127 downto 0);
signal instrs : sig_array := (
X"ca708093dff101132ef1819300000000",
X"f3a20213694282930003031300000001",
X"a6238393fff40413c2b4849300000001",
X"0ac5051345858593fff6061300000001",
X"00168693022707131827879300000001",
X"41080813912888939669091300000001",
X"3e298993fffa0a132a0a8a9300000001",
X"ff7b0b13f59b8b93d7fc0c1300000001",
X"006c8c93effd0d13d15d8d9300000001",
X"d3ee0e1386ee8e93223f0f1300000001",
X"d93f8f93000000130000001300000001",
X"00000013000000130000001300000001",
X"02c00d6f000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e0000007e0000007efffffff2"
);

type sig_array_beq_nottake is array (1 to 18) of std_logic_vector(127 downto 0);
signal instrs_beq_nottake : sig_array_beq_nottake := (
X"9eb08093842101138071819300000000",
X"f7120213de8282932a83031300000001",
X"a413839304040413acc4849300000001",
X"64750513000585933576061300000001",
X"0006869320a707136187879300000001",
X"08380813b8b88893ffd9091300000001",
X"fff98993c7fa0a13052a8a9300000001",
X"cf7b0b13dfcb8b93fefc0c1300000001",
X"311c8c937f7d0d13359d8d9300000001",
X"000e0e13551e8e93ab8f0f1300000001",
X"885f8f93000000130000001300000001",
X"00000013000000130000001300000001",
X"031b0463000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e0000007e0000007efffffff2"
);

type sig_array_beq_take is array (1 to 18) of std_logic_vector(127 downto 0);
signal instrs_beq_take : sig_array_beq_take := (
X"000080938a2101130001819300000000",
X"fef20213fff2829300a3031300000001",
X"bff38393809404130044849300000001",
X"4005051300058593a2e6061300000001",
X"06a68693fff707131d37879300000001",
X"de380813f558889305c9091300000001",
X"bf7989936b0a0a13190a8a9300000001",
X"073b0b13deab8b93040c0c1300000001",
X"fffc8c93fffd0d13fffd8d9300000001",
X"fffe0e13d92e8e93a00f0f1300000001",
X"d5ff8f93000000130000001300000001",
X"00000013000000130000001300000001",
X"02e70463000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e0000007e0000007efffffff2"
);

type sig_array_jalr2 is array (1 to 75) of std_logic_vector(127 downto 0);
type sig_array_jalr is array (1 to 84) of std_logic_vector(127 downto 0);
type sig_array_lw is array (1 to 13) of std_logic_vector(127 downto 0);

signal instrs_jalr : sig_array_jalr := (
X"ffff80b7a2410113bd11819300000000",
X"b0020213495282930e13031300000001",
X"88838393766404130004849300000001",
X"00050513082585930006061300000001",
X"df768693e9d70713df77879300000001",
X"8f38081344188893fff9091300000001",
X"88098993bfba0a13f5fa8a9300000001",
X"000b0b138cfb8b93f50c0c1300000001",
X"fffc8c936fed0d131a0d8d9300000001",
X"bbbe0e131bbe8e930a1f0f1300000001",
X"ffff8f93000000130000001300000001",
X"00000013000000130000001300000001",
X"3c808de7000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e0000007e0000007efffffff2"
);

signal instrs_jalr2 : sig_array_jalr2 := (
X"020080939a8101134dc1819300000000",
X"edf2021316e28293fbf3031300000001",
X"3c538393e7d404134814849300000001",
X"d5b50513000585931006061300000001",
X"04468693ffb707134087879300000001",
X"bff8081330088893ac79091300000001",
X"7bf98993000a0a13fdba8a9300000001",
X"fefb0b13f9db8b93504c0c1300000001",
X"004c8c93ddfd0d13fffd8d9300000001",
X"fbfe0e13dffe8e93040f0f1300000001",
X"ffaf8f93000000130000001300000001",
X"00000013000000130000001300000001",
X"36400a67000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e0000007e0000007efffffff2"
);


signal instrs_lw : sig_array_lw := (
X"4080049300000013000013b700000000",
X"82838393f277f0b77d30809300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"0093a023000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130003a08300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"00000013000000130000001300000001",
X"0000007e0000007e0000007efffffff2"
);

begin

  DUT: entity work.CPU_Comp
  generic map(N_SENSORS => 5)
  port map ( 
    system_clk            => clk,
    timer_clk             => '1',
    reset_n               => reset_n,
    
    Din                   => Din,  -- sim
    Drdy                  => Drdy, -- sim
    bsy                   => bsy,
    fsm_dvld              => fsm_dvld,
    dvld_mux              => dvld_mux,
    sensor_fifo_dvld      => sensor_fifo_dvld, -- sim

    input_data            => Kin, -- sim
    krdy                  => krdy, -- sim
    kvld                  => kvld,

    calib_trg             => calib_trg,
    sens_calib_id         => sens_calib_id,
    sensor_fifo_read      => sensor_fifo_read,
    sensor_trigger        => sensor_trigger,
    osc_trigger           => osc_trigger,
    reset_fifo            => reset_fifo,

    instruction_processed => instruction_processed,
    en_cpu                => en_cpu 

  );
        
  clk_gen: process
  begin
    clk <= '1', '0' after 50 ns;
    wait for 100 ns;
  end process;

  tb : PROCESS
  BEGIN

    reset_n <= '0';
    Kin <= (others => '0');
    Din <= (others => '0');
    Drdy <= '0';
    krdy <= '0';
    sensor_fifo_dvld <= '0';
    
    wait for 620 ns;
    
    reset_n <= '1';
    
    wait for 1000 ns;
    
    for calib in 1 to 5 loop
      -- calibration
      Kin <= X"00000000000000000000000000000003";
      krdy <= '1';
      wait for 100 ns;
      krdy <= '0';
      
      wait for 1000 ns;
      
      -- set IDC_IDF
      Kin <= X"fff000000000000000000000fffff000";
      krdy <= '1';
      wait for 100 ns;
      krdy <= '0';
      
      wait for 10000 ns;
      
      -- read a couple of sensor traces
      for i in 0 to 5 loop
        Din <= X"fffffffffffffffffffffffffffffffe";
        Drdy <= '1';
        wait for 100 ns;
        Drdy <= '0';
        
        wait until sensor_fifo_read = '1';
        wait for 500 ns;
        sensor_fifo_dvld <= '1';
        wait for 100 ns;
        sensor_fifo_dvld <= '0';
        
        wait for 1000 ns;
      end loop;
    
      -- end read of sensor traces
      Din <= X"ffffffffffffffffffffffffffffffff";
      Drdy <= '1';
      wait for 100 ns;
      Drdy <= '0';
      
      wait until dvld_mux = '1';
      
      wait for 1000 ns;
    
    end loop;
    
    wait for 10000 ns;
    
    -- rst CPU
    Kin <= X"00000000000000000000000000000007";
    krdy <= '1';
    wait for 100 ns;
    krdy <= '0';
    
    wait for 30000 ns;
    
    -- send instructions
    for i in 1 to 18 loop

        Kin <= instrs_beq_take(i);
        krdy <= '1';
        wait for 100 ns;
        krdy <= '0';
        
        wait for 1000 ns;
    end loop;
    
    Kin <= X"0000007e0000007e0000007efffffff2";
    krdy <= '1';
    wait for 100 ns;
    krdy <= '0';
    
    wait for 20000 ns;
    
    -- Offset FIFO
    --Din <= X"fffffffffffffffffffffffffff00afc";
    Din <= X"fffffffffffffffffffffffffff03ffc";
    Drdy <= '1';
    wait for 100 ns;
    Drdy <= '0';
    
    for i in 0 to 62 loop
      wait until sensor_fifo_read = '1';
      wait for 500 ns;
      sensor_fifo_dvld <= '1';
      wait for 100 ns;
      sensor_fifo_dvld <= '0';     
    end loop;
    
    wait for 20000 ns;
    
    -- Read rest of sensor traces
    for i in 0 to 5 loop
        Din <= X"fffffffffffffffffffffffffffffffe";
        Drdy <= '1';
        wait for 100 ns;
        Drdy <= '0';
        
        wait until sensor_fifo_read = '1';
        wait for 500 ns;
        sensor_fifo_dvld <= '1';
        wait for 100 ns;
        sensor_fifo_dvld <= '0';
        
        wait for 1000 ns;
    end loop;
    
    Din <= X"ffffffffffffffffffffffffffffffff";
    Drdy <= '1';
    wait for 100 ns;
    Drdy <= '0';
    
    wait until dvld_mux = '1';
    
    wait for 10000 ns;

    wait for 10000 ns;
    
    -- rst CPU
    Kin <= X"00000000000000000000000000000007";
    krdy <= '1';
    wait for 100 ns;
    krdy <= '0';
    
    wait for 30000 ns;
    
    -- send instructions
    for i in 1 to 18 loop

        Kin <= instrs_beq_take(i);
        krdy <= '1';
        wait for 100 ns;
        krdy <= '0';
        
        wait for 1000 ns;
    end loop;
    
    Kin <= X"0000007e0000007e0000007efffffff2";
    krdy <= '1';
    wait for 100 ns;
    krdy <= '0';
    
    wait for 20000 ns;
    
    -- Offset FIFO
    --Din <= X"fffffffffffffffffffffffffff00afc";
    Din <= X"fffffffffffffffffffffffffff03ffc";
    Drdy <= '1';
    wait for 100 ns;
    Drdy <= '0';
    
    for i in 0 to 62 loop
      wait until sensor_fifo_read = '1';
      wait for 500 ns;
      sensor_fifo_dvld <= '1';
      wait for 100 ns;
      sensor_fifo_dvld <= '0';     
    end loop;
    
    wait for 20000 ns;
    
    -- Read rest of sensor traces
    for i in 0 to 5 loop
        Din <= X"fffffffffffffffffffffffffffffffe";
        Drdy <= '1';
        wait for 100 ns;
        Drdy <= '0';
        
        wait until sensor_fifo_read = '1';
        wait for 500 ns;
        sensor_fifo_dvld <= '1';
        wait for 100 ns;
        sensor_fifo_dvld <= '0';
        
        wait for 1000 ns;
    end loop;
    
    Din <= X"ffffffffffffffffffffffffffffffff";
    Drdy <= '1';
    wait for 100 ns;
    Drdy <= '0';
    
    wait until dvld_mux = '1';
    
    wait for 10000 ns;
    

    wait; -- will wait forever
  END PROCESS tb;


end Behavioral;
